`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    12:46:46 04/23/2013 
// Design Name: 
// Module Name:    sprite 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module sprite( sprite, addr
    );
	 
	 input [3:0] addr;
	 output [0:31] sprite;
	 
	 reg [0:31] rom[15:0];
	 
	 initial
		begin
		
			rom[0] = 32'b01111110000011000001101000000010;
			rom[1] = 32'b01000001000011000001101000000010;
			rom[2] = 32'b01000000100010100010101000000010;
			rom[3] = 32'b01000000010010100010101000000010;
			rom[4] = 32'b01000000001010100010101000000010;
			rom[5] = 32'b01000000001010010100101000000010;
			rom[6] = 32'b01000000001010010100101000000010;
			rom[7] = 32'b01000000001010010100101111111110;
			rom[8] = 32'b01000000001010001000101000000010;
			rom[9] = 32'b01000000001010001000101000000010;
			rom[10] = 32'b01000000001010001000101000000010;
			rom[11] = 32'b01000000001010001000101000000010;
			rom[12] = 32'b01000000010010000000101000000010;
			rom[13] = 32'b01000000100010000000101000000010;
			rom[14] = 32'b01000001000010000000101000000010;
			rom[15] = 32'b01111110000010000000101000000010;
		
		end
		
	assign sprite = rom[addr];


endmodule
